`timescale 1ns / 1ps


module anodeControl(
    output reg [3:0] anode = 0,
    input [1:0] refreshCounter
    );
    
    always@(refreshCounter)
    begin
        case(refreshCounter)
            2'b00:
                anode = 4'b0111;
            2'b01:
                anode = 4'b1011;
            2'b10:
                anode = 4'b1101;
            2'b11:
                anode = 4'b1110;
        endcase
    end
endmodule